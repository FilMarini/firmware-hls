../../..//IntegrationTests/common/hdl/tf_lut.vhd