../../..//IntegrationTests/common/hdl/FileWriterFromRAM.vhd