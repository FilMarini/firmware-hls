../../..//IntegrationTests/common/hdl/FileReader.vhd