../../..//IntegrationTests/common/hdl/FileWriterFromRAMBinned.vhd