../../..//IntegrationTests/common/hdl/latency_monitor.vhd