../../..//IntegrationTests/common/hdl/FileWriter.vhd