../../..//IntegrationTests/common/hdl/tf_mem_bin.vhd