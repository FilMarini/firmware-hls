../../..//IntegrationTests/common/hdl/CreateStartSignal.vhd