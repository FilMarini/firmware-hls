../../..//IntegrationTests/common/hdl/FileReaderFIFO.vhd