../../..//IntegrationTests/common/hdl/FileWriterFIFO.vhd