../../..//IntegrationTests/common/hdl/tf_pkg.vhd