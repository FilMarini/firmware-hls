../../..//IntegrationTests/common/hdl/tf_mem.vhd